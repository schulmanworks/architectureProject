module Instruction_Memory (
                          input [31:0] PC,
                          output reg [31:0] inst);
  always @ (PC)
    case(PC)
      // I-type instructions
      0: inst =  32'h34090005; // ori $t1, $0, 0x5
      4: inst =  32'h340a0005; // ori $t2, $0, 0x5
      8: inst =  32'h340b0008; // ori $t3, $0, 0x8
      12: inst =  32'h340c000f; // ori $t4, $0, 0xf

      // R-type
      16: inst = 32'h01496024; // and $t4, $t2, $t1
      20: inst = 32'h014b6821; // addu $t5, $t2, $t3

      // More I type but stores
      24: inst = 32'hada90000; // sw $t1, 0($t5)
      28: inst = 32'hadab0004; // sw $t3, 4($t5)

      // More I type but load
      32: inst = 32'h8daa0000; // lw $t2, 0($t5)
      36: inst = 32'h8dac0004; // lw $t4, 4($t5)
      // 0: inst =   32'b00111100000000011111111111111111; //1. lui $1, 1
      // 4: inst =   32'b00000000000000010001010000000011; //2. sra $2, $1, 16
      // 8: inst =   32'b00000000000000100001110000000000; //3. sll $3, $2, 16
      // 12: inst =  32'b00000000000000110010011000000010; //4. srl $4, $3, 24
      // 16: inst =  32'b00100100000001010000000000001111; //5. addui $5, $0, 17
      // 20: inst =  32'b00000000100001010011000000100011; //6.  subu $6, $4, $5
      // 24: inst =  32'b00000000110001000011100000100001; //7.  addu $7, $6, $4
      // 28: inst =  32'b00000000111001100100000000100100; //8.  and  $8, $7, $6
      // 32: inst =  32'b00000000111001100100100000100110; //9.  xor  $9, $7, $6
      // 36: inst =  32'b00000000001010010101000000101010; //10. slt  $10, $1, $9
      // 40: inst =  32'b00010101010000000000000000000010; //11. bne  $10, $0, xxx,
      // // next instruction is 52 = PC+4 + 8
      //
      // 52: inst =  32'b00000000111010010101100000100101; //12  or  $11, $7, $9
      // 56: inst =  32'b00001100000000000000000000010010; //13  jal XXXX
      // // I'll jump C0 72 = 1001000
      // 72: inst =  32'b00110001011011000000000000001010; //14. andi $12, $11, 1010
      // 76: inst =  32'b00000011111000000000000000001000; //15. jr $31
      // // next instruction is 60 [56+4: inst from $31
      // 60: inst =  32'b00001000000000000000000000010100; //16. j zzzz
      // // next instruction is 80 = 1010000
      // 80: inst =  32'b10001101100011010000000000000000; //17. lw  $13, 0($12)
      // 84: inst =  32'b00111001101011100000000000001110; //18. xori $14, $13, 1110
      // 88: inst =  32'b00110101101011110000000000001110; //19. ori  $15, $13, 1110
      // 92: inst =  32'b00000000001010011000000000101011; //20. sltu $16, $1, $9
      // 96: inst =  32'b00101000001100010000000000000000; //21. slti $17, $1, 0
      // 100: inst = 32'b00101100001100100000000000000000; //22. sltui $18, s1, 0
      // 104: inst = 32'b00010010000100100000000000000010; //23. beq $16,$18, yyyy
      // // next instruction is +12 (4+8)
      // 116: inst = 32'b10101101100010110000000000000100; //24. sw $11, 4(12)
      default: inst = 32'b0;
    endcase
endmodule
